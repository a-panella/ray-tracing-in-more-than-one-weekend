context rt_sim_context is
    library rt;
    context rt.rt_context;
    use rt.sim_pkg.all;
    library ieee;
    use std.textio.all;
    -- include OSVVM packages here when using them later...
end context;