context rt_context is
    library rt;
    context rt.rt_base_context;
    use rt.src_pkg.all;
end context;

